library verilog;
use verilog.vl_types.all;
entity arf_vlg_vec_tst is
end arf_vlg_vec_tst;
